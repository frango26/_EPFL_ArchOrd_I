library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity register_file is
	port(
		clk    : in std_logic;
		aa     : in  std_logic_vector( 4 downto 0);
		ab     : in  std_logic_vector( 4 downto 0);
		aw     : in  std_logic_vector( 4 downto 0);
		wren   : in  std_logic;
		wrdata : in  std_logic_vector(31 downto 0);
		a      : out std_logic_vector(31 downto 0);
		b      : out std_logic_vector(31 downto 0)
	);
end register_file;

architecture synth of register_file is
begin
	
end synth;
