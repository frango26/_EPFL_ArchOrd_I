library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity add_sub is
	port(
		a        : in  std_logic_vector(31 downto 0);
		b        : in  std_logic_vector(31 downto 0);
		sub_mode : in  std_logic;
		carry    : out std_logic;
		zero     : out std_logic;
		r        : out std_logic_vector(31 downto 0)
	);
end add_sub;

architecture synth of add_sub is

begin

end synth;