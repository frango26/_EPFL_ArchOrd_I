library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity comparator is
	port (
		a_31    : in  std_logic;
		b_31    : in  std_logic;
		diff_31 : in  std_logic;
		carry   : in  std_logic;
		zero    : in  std_logic;
		op      : in  std_logic_vector( 2 downto 0);
		r       : out std_logic
	);
end comparator;

architecture synth of comparator is

begin

end synth;
