library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity ROM is
	port(
		clk     : in  std_logic;
		cs      : in  std_logic;
		read    : in  std_logic;
		address : in  std_logic_vector(9 downto 0);
		rddata  : out std_logic_vector(31 downto 0));
end ROM;

architecture synth of ROM is
begin
	rddata <= (others => 'Z');
end synth;
